(* TODO: rename to LLVMCFG? *)
Require Import Equalities.

From Coq Require Import ZArith List String.

From SE Require Import
     Utilities
     LLVMAst.

From ExtLib Require Import
     Programming.Eqv
     Structures.Monads.

Import ListNotations.
Import EqvNotation.
Import MonadNotation.
Open Scope list.
Open Scope monad_scope.

Section CFG.

  Variable (T:Set).

  Record cfg := mk_cfg {
    init : block_id;
    blks : list (block T);
  }.

  Record module {Body : Set} : Set := mk_module {
    m_name : option string;
    m_target : option string;
    m_datalayout : option string;
    m_type_defs : list (ident * T);
    m_globals : list (global T);
    m_declarations : list (declaration T);
    m_definitions : list (@definition T Body);
  }.

End CFG.

Arguments mk_cfg {_}.
Arguments init {_}.
Arguments blks {_}.
Arguments module {_} _.
Arguments mk_module {_ _}.
Arguments m_name {_ _}.
Arguments m_target {_ _}.
Arguments m_datalayout {_ _}.
Arguments m_type_defs {_ _}.
Arguments m_globals {_ _}.
Arguments m_declarations {_ _}.
Arguments m_definitions {_ _}.

Definition llvm_exp := @exp typ.
Definition llvm_global := @global typ.
Definition llvm_cmd := @cmd typ.
Definition llvm_block := @block typ.
Definition llvm_cfg := @cfg typ.
Definition llvm_declaration := @declaration typ.
Definition llvm_definition := @definition typ llvm_cfg.
Definition llvm_module : Set := @module typ llvm_cfg.

Definition get_cmd_id (c : llvm_cmd) : cmd_id :=
  match c with
  | CMD_Phi n _ => n
  | CMD_Inst n _ => n
  | CMD_Term n _ => n
  end
.

Definition get_first_cmd (b : llvm_block) : option cmd :=
  match (blk_cmds b) with
  | c :: _ => Some c
  | _ => None
  end
.

Definition get_first_cmd_id (b : llvm_block) : option cmd_id :=
  match (get_first_cmd b) with
  | Some c => Some (get_cmd_id c)
  | _ => None
  end
.

Definition match_block (bid : block_id) (b : llvm_block) : bool :=
  if (blk_id b) =? bid then true else false
.

Definition find_block (bs: list (llvm_block)) (bid : block_id) : option (llvm_block) :=
  find (fun b => match_block bid b) bs
.

(* TODO: rename *)
Definition get_fid(d : llvm_definition) : function_id :=
  (dc_name (df_prototype d))
.

Definition fetch_block (d : llvm_definition) (bid : block_id) : option llvm_block :=
  find_block (blks (df_body d)) bid
.

Definition entry_block (d : llvm_definition) : option llvm_block :=
  fetch_block d (init (df_body d))
.

Definition match_declaration (fid : function_id) (d : llvm_declaration) : option (llvm_declaration) :=
  if (dc_name d) =? fid then Some d else None
.

Definition find_declaration (m : llvm_module) (fid : function_id) : option (llvm_declaration) :=
  find_map (match_declaration fid) (m_declarations m)
.

Definition match_function (fid : function_id) (d : llvm_definition) : option (llvm_definition) :=
  if (dc_name (df_prototype d)) =? fid then Some d else None
.

Definition find_function (m : llvm_module) (fid : function_id) : option (llvm_definition) :=
  find_map (match_function fid) (m_definitions m)
.

Definition find_function_by_exp (m : llvm_module) (e : llvm_exp) : option llvm_definition :=
  match e with
  | EXP_Ident (ID_Global id) => find_function m id
  | _ => None
  end
.

(* TODO: rename *)
Lemma LX1 : forall mdl d fid,
  find_function mdl fid = Some d ->
  In d (m_definitions mdl).
Proof.
Admitted.

(* TODO: rename *)
Lemma LX2 : forall d bid b,
  fetch_block d bid = Some b ->
  In b (blks (df_body d)).
Proof.
Admitted.

Inductive llvm_subexpr : llvm_exp -> llvm_exp -> Prop :=
  | LLVM_SubExpr_Refl : forall e, llvm_subexpr e e
  | LLVM_SubExpr_Trans : forall e1 e2 e3,
      llvm_subexpr e1 e2 -> llvm_subexpr e2 e3 -> llvm_subexpr e1 e3
  | LLVM_SubExpr_IBinop_L : forall op t e1 e2,
      llvm_subexpr e1 (OP_IBinop op t e1 e2)
  | LLVM_SubExpr_IBinop_R : forall op t e1 e2,
      llvm_subexpr e2 (OP_IBinop op t e1 e2)
  | LLVM_SubExpr_ICmp_L : forall op t e1 e2,
      llvm_subexpr e1 (OP_ICmp op t e1 e2)
  | LLVM_SubExpr_ICmp_R : forall op t e1 e2,
      llvm_subexpr e2 (OP_ICmp op t e1 e2)
  | LLVM_SubExpr_Conversion : forall conv t1 t2 e,
      llvm_subexpr e (OP_Conversion conv t1 e t2)
  | LLVM_SubExpr_Select_Cond : forall t1 e1 t2 e2 t3 e3,
      llvm_subexpr e1 (OP_Select (t1, e1) (t2, e2) (t3, e3))
  | LLVM_SubExpr_Select_L : forall t1 e1 t2 e2 t3 e3,
      llvm_subexpr e2 (OP_Select (t1, e1) (t2, e2) (t3, e3))
  | LLVM_SubExpr_Select_R : forall t1 e1 t2 e2 t3 e3,
      llvm_subexpr e3 (OP_Select (t1, e1) (t2, e2) (t3, e3))
.
